module ysyx_25040129_MMU (
	input clk,
	input rst,
	input [31:0] satp

	
);
	
endmodule