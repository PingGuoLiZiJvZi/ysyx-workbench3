module ysyx_25040129_UART(

);

endmodule
